* source INV
M_M1         OUT N14434 0 0 NMOS  
+ L=.18u  
+ W=.76u         
M_M2         OUT N14434 N14461 N14461 PMOS  
+ L=.18u  
+ W=1.8u         
V_V1         N14461 0 1.8Vdc
V_V2         N14434 0  
+PULSE 1.8V 0V 0ns 1ns 1ns 2us 4us
C_C1         0 OUT  20p 
.MODEL PMOS PMOS
.MODEL NMOS NMOS  
.tran 2e-0 20e-6 2e-6 
.control
run
plot V(out) 
.endc
.end