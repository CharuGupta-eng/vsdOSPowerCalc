* source MUX
M_M5         A SEL OUT VDD Mbreakp  
+ L=.18u  
+ W=1.8u         
M_M4         OUT SEL B 0 Mbreakn  
+ L=.18u  
+ W=.72u         
V_V6         SEL 0  
+PULSE 1.8V 0 0 1n 1n 1u 2u
V_V10         A 0  
+PULSE 1.8V 0V 0 1n 1n 3u 6u
V_V11         B 0  
+PULSE 1.8V 0V 0 1n 1n 2u 4u
V_V5         VDD 0 1.8Vdc
C_C2         0 OUT  20p  

.MODEL MBREAKP PMOS
.MODEL MBREAKN NMOS  
.tran 2e-0 20e-6 
.control
run 
PLOT V(OUT)
PLOT V(SEL)
PLOT V(A)
PLOT V(B)

.endc
.end 
