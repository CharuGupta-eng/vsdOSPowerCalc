* source NET_DFF_PT
V_V17         DIN 0  
M_M13         N40957 N40799 VDD VDD MbreakP  
+ L=.18u  
+ W=.72u         
M_M14         QBAR N41061 0 0 MbreakN  
+ L=.18u  
+ W=.72u         
M_M10         N40799 N40739 0 0 Mbreakn  
+ L=.18u  
+ W=.72u         
M_M18         N40739 CLK DIN 0 MbreakN  
+ L=.18u  
+ W=.72u         
M_M16         Q QBAR 0 0 MbreakN  
+ L=.18u  
+ W=.72u         
M_M15         QBAR N41061 VDD VDD MbreakP  
+ L=.18u  
+ W=.72u         
M_M19         N40957 CLK N40739 VDD MbreakP  
+ L=.18u  
+ W=.72u         
M_M12         N40957 N40799 0 0 MbreakN  
+ L=.18u  
+ W=.72u         
M_M20         Q CLK N41061 0 MbreakN  
+ L=.18u  
+ W=.72u         
M_M17         Q QBAR VDD VDD MbreakP  
+ L=.18u  
+ W=.72u         
C_C5         0 Q  20p 
V_V18         CLK 0  
M_M11         N40799 N40739 VDD VDD Mbreakp  
+ L=.18u  
+ W=.72u         
M_M21         N41061 CLK N40957 VDD MbreakP  
+ L=.18u  
+ W=.72u         
V_V12         N43383 0 1.8Vdc
V_V19         N43383 VDD 0Vdc
   
.MODEL MBREAKP PMOS
.MODEL MBREAKN NMOS  
.OP
.control
run 
PLOT V(Q)
PLOT V(CLK)
PLOT V(DIN)
PLOT V(VDD)* I(V_V19)
PRINT V(VDD)* I(V_V19)
.endc
.end  