* source MUX_TG
M_M8         OUTPUTTG N22714 B VDD MbreakP  
+ L=.18u  
+ W=.72u         
C_C2         0 OUTPUTTG  20p  
M_M5         N22714 SEL N22696 N22696 Mbreakp  
+ L=.18u  
+ W=1.8u         
M_M4         N22714 SEL 0 0 Mbreakn  
+ L=.18u  
+ W=.72u         
V_V6         SEL 0  
M_M7         A N22714 OUTPUTTG 0 MbreakN  
+ L=.18u  
+ W=.72u         
V_V10         A 0  
V_V11         B 0  
M_M9         B SEL OUTPUTTG 0 MbreakN  
+ L=.18u  
+ W=.72u         
M_M6         OUTPUTTG SEL A VDD MbreakP  
+ L=.18u  
+ W=.72u         
V_V5         N24354 0 1.8Vdc
V_V12         N24354 VDD 0Vdc      
.MODEL MBREAKP PMOS
.MODEL MBREAKN NMOS  
.op
.control
run 
PLOT V(OUTPUTTG)
PLOT V(SEL)
PLOT V(A)
PLOT V(B)
PLOT V(VDD)* I(V_V12)
PRINT V(VDD)* I(V_V12)
.endc
.end  