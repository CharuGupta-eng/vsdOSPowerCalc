* source INV
M_M1         OUT N14434 0 0 NMOS  
+ L=.18u  
+ W=.76u         
M_M2         OUT N14434 VD VD PMOS  
+ L=.18u  
+ W=1.8u         
V_V1         VDD 0 1.8Vdc
V_V2         N14434 0  
C_C1         0 OUT  20p   
V_V3         VDD VD 0Vdc
   
.MODEL PMOS PMOS
.MODEL NMOS NMOS  
.op
.control
run
plot V(out)
plot V(VDD)
print I(V_V3)* V(VDD) 
.endc
.end