10bitdac
V1 N001 0 3.3
XX1 d0 d1 d2 d3 d4 d5 d6 d7 d8 d9 out N002 0 level9
R1 N001 N002 5k
V2 d0 0 0
V3 d1 0 0
V4 d2 0 0
V5 d3 0 0
V6 d4 0 0
V7 d5 0 0
V8 d6 0 0
V9 d7 0 0
V10 d8 0 0
V11 d9 0 0

* block symbol definitions
.subckt level9 d0 d1 d2 d3 d4 d5 d6 d7 d8 d9 out_10 res_in10 res_out10
XX1 d0 d1 d2 d3 d4 d5 d6 d7 d8 res_in10 N002 N001 level8
XX2 d0 d1 d2 d3 d4 d5 d6 d7 d8 N003 res_out10 N004 level8
XX3 d9 N001 N004 out_10 switch
R1 N002 N003 5k
.ends level9

.subckt level8 d0 d1 d2 d3 d4 d5 d6 d7 d8 res_in9 res_out9 out_9
XX1 d0 d1 d2 d3 d4 d5 d6 d7 N002 N001 res_in9 level7
XX2 d0 d1 d2 d3 d4 d5 d6 d7 res_out9 N004 N003 level7
XX3 d8 N001 N004 out_9 switch
R1 N002 N003 5k
.ends level8

.subckt switch dig_in in_1 in_2 Vout
M1 in_1 dig_in Vout Vout CMOSN L=180n W =360n
M2 Vout N002 in_2 in_2 CMOSN L=180n W =360n
M4 N002 dig_in 0 0 CMOSN L=180n W =360n
M5 N002 dig_in N001 N001 CMOSP L=180n W =900n
M6 in_2 dig_in Vout Vout CMOSP L=180n W =900n
M3 Vout N002 in_1 in_1 CMOSP L=180n W =900n
V1 N001 0 3.3
.model CMOSN NMOS (LEVEL=8 VERSION=3.2 TNOM=27 TOX=4.1E-9 XJ=1E-7 NCH=2.3549E17 VTH0=0.3823463 K1=0.5810697 
+            K2=4.774618E-3 K3=0.0431669 K3B=1.1498346 W0=1E-7 NLX=1.910552E-7 DVT0W=0 DVT1W=0 DVT2W=0 
+            DVT0=1.2894824 DVT1=0.3622063 DVT2=0.0713729 U0=280.633249 UA=-1.208537E-9 UB=2.158625E-18
+            UC=5.342807E-11 VSAT=9.366802E4 A0=1.7593146 AGS=0.3939741 B0=-6.413949E-9 B1=-1E-7 KETA=-5.180424E-4
+            A1=0 A2=1 RDSW=105.5517558 PRWG=0.5 PRWB=-0.1998871 WR=1 WINT=7.904732E-10 LINT=1.571424E-8 XL=0
+            XW=-1E-8 DWG=1.297221E-9 DWB=1.479041E-9 VOFF=-0.0955434 NFACTOR=2.4358891 CIT=0 CDSC=2.4E-4 CDSCD=0
+            CDSCB=0 ETA0=3.104851E-3 ETAB=-2.512384E-5 DSUB=0.0167075 PCLM=0.8073191 PDIBLC1=0.1666161 PDIBLC2=3.112892E-3    
+            PDIBLCB=-0.1 DROUT=0.7875618 PSCBE1=8E10 PSCBE2=9.213635E-10 PVAG=3.85243E-3 DELTA=0.01 RSH=6.7 MOBMOD=1
+            PRT=0 UTE=-1.5 KT1=-0.11 KT1L=0 KT2=0.022 UA1=4.31E-9 UB1=-7.61E-18 UC1=-5.6E-11 AT=3.3E4 WL=0 WLN=1
+            WW=0 WWN=1 WWL=0 LL=0 LLN=1 LW=0 LWN=1 LWL=0 CAPMOD=2 XPART=0.5 CGDO=7.08E-10 CGSO=7.08E-10 CGBO=1E-12
+            CJ=9.68858E-4 PB=0.8 MJ=0.3864502 CJSW=2.512138E-10 PBSW=0.809286 MJSW=0.1060414 CJSWG=3.3E-10 PBSWG=0.809286 
+            MJSWG=0.1060414 CF=0 PVTH0=-1.192722E-3 PRDSW=-5 PK2=6.450505E-5 WKETA=-4.27294E-4 LKETA=-0.0104078 
+            PU0=6.3268729 PUA=2.226552E-11 PUB=0 PVSAT=969.1480157 PETA0=1E-4 PKETA=-1.049509E-3)

.model CMOSP PMOS (LEVEL=8 VERSION=3.2 TNOM=27 TOX=4.1E-9 XJ=1E-7 NCH=4.1589E17 VTH0=-0.3938813 K1=0.5479015
+            K2=0.0360586 K3=0.0993095 K3B=5.7086622 W0=1E-6 NLX=1.313191E-7 DVT0W=0 DVT1W=0 DVT2W=0 DVT0=0.4911363
+            DVT1=0.2227356 DVT2=0.1 U0=115.6852975 UA=1.505832E-9 UB=1E-21 UC=-1E-10 VSAT=1.329694E5 A0=1.7590478
+            AGS=0.3641621 B0=3.427126E-7 B1=1.062928E-6 KETA=0.0134667 A1=0.6859506 A2=0.3506788 RDSW=168.5705677
+            PRWG=0.5 PRWB=-0.4987371 WR=1 WINT=0 LINT=3.028832E-8 XL=0 XW=-1E-8 DWG=-2.349633E-8 DWB=-7.152486E-9 
+            VOFF=-0.0994037 NFACTOR=1.9424315 CIT=0 CDSC=2.4E-4 CDSCD=0 CDSCB=0 ETA0=0.0608072 ETAB=-0.0426148
+            DSUB=0.7343015 PCLM=3.2579974 PDIBLC1=7.229527E-6 PDIBLC2=0.025389 PDIBLCB=-1E-3 DROUT=0 PSCBE1=1.454878E10
+            PSCBE2=4.202027E-9 PVAG=15 DELTA=0.01 RSH=7.8 MOBMOD=1 PRT=0 UTE=-1.5 KT1=-0.11 KT1L=0 KT2=0.022 UA1=4.31E-9
+            UB1=-7.61E-18 UC1=-5.6E-11 AT=3.3E4 WL=0 WLN=1 WW=0 WWN=1 WWL=0 LL=0 LLN=1 LW=0 LWN=1 LWL=0 CAPMOD=2 XPART=0.5
+            CGDO=6.32E-10 CGSO=6.32E-10 CGBO=1E-12 CJ=1.172138E-3 PB=0.8421173 MJ=0.4109788 CJSW=2.242609E-10 PBSW=0.8            
+            MJSW=0.3752089 CJSWG=4.22E-10 PBSWG=0.8 MJSWG=0.3752089 CF=0 PVTH0=1.888482E-3 PRDSW=11.5315407 PK2=1.559399E-3    
+            WKETA=0.0319301 LKETA=2.955547E-3 PU0=-1.1105313 PUA=-4.62102E-11 PUB=1E-21 PVSAT=50 PETA0=1E-4 PKETA=-4.346368E-3)

.ends switch

.subckt level7 d0 d1 d2 d3 d4 d5 d6 d7 res_out8 out_8 res_in8
XX1 d0 d1 d2 d3 d4 d5 d6 res_in8 N002 N001 level6
XX2 d0 d1 d2 d3 d4 d5 d6 N003 res_out8 N004 level6
XX3 d7 N001 N004 out_8 switch
R1 N002 N003 5k
.ends level7

.subckt level6 d0 d1 d2 d3 d4 d5 d6 res_in7 res_out7 out_7
XX1 d0 d1 d2 d3 d4 d5 res_in7 N002 N001 level5
XX2 d0 d1 d2 d3 d4 d5 N003 res_out7 N004 level5
R1 N002 N003 5k
XX3 d6 N001 N004 out_7 switch
.ends level6

.subckt level5 d0 d1 d2 d3 d4 d5 res_in6 res_out6 out_6
XX1 d0 d1 d2 d3 d4 res_in6 N002 N001 level4
XX2 d0 d1 d2 d3 d4 N003 res_out6 N004 level4
XX3 d5 N001 N004 out_6 switch
R1 N002 N003 5k
.ends level5

.subckt level4 d0 d1 d2 d3 d4 str_in str_out out_5
XX1 d0 d1 d2 d3 str_in P001 N001 level3
XX2 d0 d1 d2 d3 N002 str_out N003 level3
XX3 d4 N001 N003 out_5 switch
R1 P001 N002 5k
.ends level4

.subckt level3 d0 d1 d2 d3 res_in res_out output
XX1 d0 d1 d2 res_in N002 N001 level2
XX2 d0 d1 d2 N003 res_out N004 level2
XX3 d3 N001 N004 output switch
R1 N002 N003 5k
.ends level3

.subckt level2 d0 d1 d2 in_res out_res out
XX1 in_res N002 N001 d0 d1 level1
XX2 N003 out_res N004 d0 d1 level1
XX3 d2 N001 N004 out switch
R1 N002 N003 5k
.ends level2

.subckt level1 in_pin out_pin out_v d0 d1
XX1 d0 in_pin N002 N001 switch
XX2 d0 N003 N005 N004 switch
XX3 d1 N001 N004 out_v switch
R1 in_pin N002 10k
R2 N005 out_pin 5k
R3 N002 N003 10k
R4 N003 N005 10k
.ends level1


.tran 100e-03 8e-00 0e-00
* Control Statements 
.control
run
plot v(out)
.endc
.end