* source NET_MUX_2T
V_V1         A 0  
+PULSE 1.8V 0 0 1n 1n 3u 6u
V_V2         SEL 0  
+PULSE 1.8V 0V 0 1n 1n 1u 2u
M_M1         OUT SEL B 0 Mbreakn  
+ L=.18u  
+ W=.72u         
M_M3         A SEL OUT VDD Mbreakp  
+ L=.18u  
+ W=.72u         
V_V4         N15973 0 1.8Vdc
V_V3         B 0  
+PULSE 1.8V 0V 0 1n 1n 2u 4u
C_C1         0 OUT  20p  
V_V5         N15973 VDD 0Vdc 
F1 0 5 V_V5 0.09
C1 5 0 10n
R1 5 0 100K  
.MODEL MBREAKP PMOS
.MODEL MBREAKN NMOS  
.tran 2e-0 20e-6 uic
.control
run 
*PLOT V(OUT)
*PLOT V(SEL)
*PLOT V(A)
*PLOT V(B)
*PLOT V(VDD) * I(V_V5)
*PRINT V(VDD) * I(V_V5)
PLOT V(5)
PRINT V(5)
.endc
.end  